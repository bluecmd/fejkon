10'b1001110100 : symbol <= "D00.0 -";
10'b0110001011 : symbol <= "D00.0 +";
10'b1001111001 : symbol <= "D00.1 -";
10'b0110001001 : symbol <= "D00.1 +";
10'b1001110101 : symbol <= "D00.2 -";
10'b0110000101 : symbol <= "D00.2 +";
10'b1001110011 : symbol <= "D00.3 -";
10'b0110001100 : symbol <= "D00.3 +";
10'b1001110010 : symbol <= "D00.4 -";
10'b0110001101 : symbol <= "D00.4 +";
10'b1001111010 : symbol <= "D00.5 -";
10'b0110001010 : symbol <= "D00.5 +";
10'b1001110110 : symbol <= "D00.6 -";
10'b0110000110 : symbol <= "D00.6 +";
10'b1001110001 : symbol <= "D00.7 -";
10'b0110001110 : symbol <= "D00.7 +";
10'b0111010100 : symbol <= "D01.0 -";
10'b1000101011 : symbol <= "D01.0 +";
10'b0111011001 : symbol <= "D01.1 -";
10'b1000101001 : symbol <= "D01.1 +";
10'b0111010101 : symbol <= "D01.2 -";
10'b1000100101 : symbol <= "D01.2 +";
10'b0111010011 : symbol <= "D01.3 -";
10'b1000101100 : symbol <= "D01.3 +";
10'b0111010010 : symbol <= "D01.4 -";
10'b1000101101 : symbol <= "D01.4 +";
10'b0111011010 : symbol <= "D01.5 -";
10'b1000101010 : symbol <= "D01.5 +";
10'b0111010110 : symbol <= "D01.6 -";
10'b1000100110 : symbol <= "D01.6 +";
10'b0111010001 : symbol <= "D01.7 -";
10'b1000101110 : symbol <= "D01.7 +";
10'b1011010100 : symbol <= "D02.0 -";
10'b0100101011 : symbol <= "D02.0 +";
10'b1011011001 : symbol <= "D02.1 -";
10'b0100101001 : symbol <= "D02.1 +";
10'b1011010101 : symbol <= "D02.2 -";
10'b0100100101 : symbol <= "D02.2 +";
10'b1011010011 : symbol <= "D02.3 -";
10'b0100101100 : symbol <= "D02.3 +";
10'b1011010010 : symbol <= "D02.4 -";
10'b0100101101 : symbol <= "D02.4 +";
10'b1011011010 : symbol <= "D02.5 -";
10'b0100101010 : symbol <= "D02.5 +";
10'b1011010110 : symbol <= "D02.6 -";
10'b0100100110 : symbol <= "D02.6 +";
10'b1011010001 : symbol <= "D02.7 -";
10'b0100101110 : symbol <= "D02.7 +";
10'b1100011011 : symbol <= "D03.0 -";
10'b1100010100 : symbol <= "D03.0 +";
10'b1100011001 : symbol <= "D03.1 -";
10'b1100011001 : symbol <= "D03.1 +";
10'b1100010101 : symbol <= "D03.2 -";
10'b1100010101 : symbol <= "D03.2 +";
10'b1100011100 : symbol <= "D03.3 -";
10'b1100010011 : symbol <= "D03.3 +";
10'b1100011101 : symbol <= "D03.4 -";
10'b1100010010 : symbol <= "D03.4 +";
10'b1100011010 : symbol <= "D03.5 -";
10'b1100011010 : symbol <= "D03.5 +";
10'b1100010110 : symbol <= "D03.6 -";
10'b1100010110 : symbol <= "D03.6 +";
10'b1100011110 : symbol <= "D03.7 -";
10'b1100010001 : symbol <= "D03.7 +";
10'b1101010100 : symbol <= "D04.0 -";
10'b0010101011 : symbol <= "D04.0 +";
10'b1101011001 : symbol <= "D04.1 -";
10'b0010101001 : symbol <= "D04.1 +";
10'b1101010101 : symbol <= "D04.2 -";
10'b0010100101 : symbol <= "D04.2 +";
10'b1101010011 : symbol <= "D04.3 -";
10'b0010101100 : symbol <= "D04.3 +";
10'b1101010010 : symbol <= "D04.4 -";
10'b0010101101 : symbol <= "D04.4 +";
10'b1101011010 : symbol <= "D04.5 -";
10'b0010101010 : symbol <= "D04.5 +";
10'b1101010110 : symbol <= "D04.6 -";
10'b0010100110 : symbol <= "D04.6 +";
10'b1101010001 : symbol <= "D04.7 -";
10'b0010101110 : symbol <= "D04.7 +";
10'b1010011011 : symbol <= "D05.0 -";
10'b1010010100 : symbol <= "D05.0 +";
10'b1010011001 : symbol <= "D05.1 -";
10'b1010011001 : symbol <= "D05.1 +";
10'b1010010101 : symbol <= "D05.2 -";
10'b1010010101 : symbol <= "D05.2 +";
10'b1010011100 : symbol <= "D05.3 -";
10'b1010010011 : symbol <= "D05.3 +";
10'b1010011101 : symbol <= "D05.4 -";
10'b1010010010 : symbol <= "D05.4 +";
10'b1010011010 : symbol <= "D05.5 -";
10'b1010011010 : symbol <= "D05.5 +";
10'b1010010110 : symbol <= "D05.6 -";
10'b1010010110 : symbol <= "D05.6 +";
10'b1010011110 : symbol <= "D05.7 -";
10'b1010010001 : symbol <= "D05.7 +";
10'b0110011011 : symbol <= "D06.0 -";
10'b0110010100 : symbol <= "D06.0 +";
10'b0110011001 : symbol <= "D06.1 -";
10'b0110011001 : symbol <= "D06.1 +";
10'b0110010101 : symbol <= "D06.2 -";
10'b0110010101 : symbol <= "D06.2 +";
10'b0110011100 : symbol <= "D06.3 -";
10'b0110010011 : symbol <= "D06.3 +";
10'b0110011101 : symbol <= "D06.4 -";
10'b0110010010 : symbol <= "D06.4 +";
10'b0110011010 : symbol <= "D06.5 -";
10'b0110011010 : symbol <= "D06.5 +";
10'b0110010110 : symbol <= "D06.6 -";
10'b0110010110 : symbol <= "D06.6 +";
10'b0110011110 : symbol <= "D06.7 -";
10'b0110010001 : symbol <= "D06.7 +";
10'b1110001011 : symbol <= "D07.0 -";
10'b0001110100 : symbol <= "D07.0 +";
10'b1110001001 : symbol <= "D07.1 -";
10'b0001111001 : symbol <= "D07.1 +";
10'b1110000101 : symbol <= "D07.2 -";
10'b0001110101 : symbol <= "D07.2 +";
10'b1110001100 : symbol <= "D07.3 -";
10'b0001110011 : symbol <= "D07.3 +";
10'b1110001101 : symbol <= "D07.4 -";
10'b0001110010 : symbol <= "D07.4 +";
10'b1110001010 : symbol <= "D07.5 -";
10'b0001111010 : symbol <= "D07.5 +";
10'b1110000110 : symbol <= "D07.6 -";
10'b0001110110 : symbol <= "D07.6 +";
10'b1110001110 : symbol <= "D07.7 -";
10'b0001110001 : symbol <= "D07.7 +";
10'b1110010100 : symbol <= "D08.0 -";
10'b0001101011 : symbol <= "D08.0 +";
10'b1110011001 : symbol <= "D08.1 -";
10'b0001101001 : symbol <= "D08.1 +";
10'b1110010101 : symbol <= "D08.2 -";
10'b0001100101 : symbol <= "D08.2 +";
10'b1110010011 : symbol <= "D08.3 -";
10'b0001101100 : symbol <= "D08.3 +";
10'b1110010010 : symbol <= "D08.4 -";
10'b0001101101 : symbol <= "D08.4 +";
10'b1110011010 : symbol <= "D08.5 -";
10'b0001101010 : symbol <= "D08.5 +";
10'b1110010110 : symbol <= "D08.6 -";
10'b0001100110 : symbol <= "D08.6 +";
10'b1110010001 : symbol <= "D08.7 -";
10'b0001101110 : symbol <= "D08.7 +";
10'b1001011011 : symbol <= "D09.0 -";
10'b1001010100 : symbol <= "D09.0 +";
10'b1001011001 : symbol <= "D09.1 -";
10'b1001011001 : symbol <= "D09.1 +";
10'b1001010101 : symbol <= "D09.2 -";
10'b1001010101 : symbol <= "D09.2 +";
10'b1001011100 : symbol <= "D09.3 -";
10'b1001010011 : symbol <= "D09.3 +";
10'b1001011101 : symbol <= "D09.4 -";
10'b1001010010 : symbol <= "D09.4 +";
10'b1001011010 : symbol <= "D09.5 -";
10'b1001011010 : symbol <= "D09.5 +";
10'b1001010110 : symbol <= "D09.6 -";
10'b1001010110 : symbol <= "D09.6 +";
10'b1001011110 : symbol <= "D09.7 -";
10'b1001010001 : symbol <= "D09.7 +";
10'b0101011011 : symbol <= "D10.0 -";
10'b0101010100 : symbol <= "D10.0 +";
10'b0101011001 : symbol <= "D10.1 -";
10'b0101011001 : symbol <= "D10.1 +";
10'b0101010101 : symbol <= "D10.2 -";
10'b0101010101 : symbol <= "D10.2 +";
10'b0101011100 : symbol <= "D10.3 -";
10'b0101010011 : symbol <= "D10.3 +";
10'b0101011101 : symbol <= "D10.4 -";
10'b0101010010 : symbol <= "D10.4 +";
10'b0101011010 : symbol <= "D10.5 -";
10'b0101011010 : symbol <= "D10.5 +";
10'b0101010110 : symbol <= "D10.6 -";
10'b0101010110 : symbol <= "D10.6 +";
10'b0101011110 : symbol <= "D10.7 -";
10'b0101010001 : symbol <= "D10.7 +";
10'b1101001011 : symbol <= "D11.0 -";
10'b1101000100 : symbol <= "D11.0 +";
10'b1101001001 : symbol <= "D11.1 -";
10'b1101001001 : symbol <= "D11.1 +";
10'b1101000101 : symbol <= "D11.2 -";
10'b1101000101 : symbol <= "D11.2 +";
10'b1101001100 : symbol <= "D11.3 -";
10'b1101000011 : symbol <= "D11.3 +";
10'b1101001101 : symbol <= "D11.4 -";
10'b1101000010 : symbol <= "D11.4 +";
10'b1101001010 : symbol <= "D11.5 -";
10'b1101001010 : symbol <= "D11.5 +";
10'b1101000110 : symbol <= "D11.6 -";
10'b1101000110 : symbol <= "D11.6 +";
10'b1101001110 : symbol <= "D11.7 -";
10'b1101001000 : symbol <= "D11.7 +";
10'b0011011011 : symbol <= "D12.0 -";
10'b0011010100 : symbol <= "D12.0 +";
10'b0011011001 : symbol <= "D12.1 -";
10'b0011011001 : symbol <= "D12.1 +";
10'b0011010101 : symbol <= "D12.2 -";
10'b0011010101 : symbol <= "D12.2 +";
10'b0011011100 : symbol <= "D12.3 -";
10'b0011010011 : symbol <= "D12.3 +";
10'b0011011101 : symbol <= "D12.4 -";
10'b0011010010 : symbol <= "D12.4 +";
10'b0011011010 : symbol <= "D12.5 -";
10'b0011011010 : symbol <= "D12.5 +";
10'b0011010110 : symbol <= "D12.6 -";
10'b0011010110 : symbol <= "D12.6 +";
10'b0011011110 : symbol <= "D12.7 -";
10'b0011010001 : symbol <= "D12.7 +";
10'b1011001011 : symbol <= "D13.0 -";
10'b1011000100 : symbol <= "D13.0 +";
10'b1011001001 : symbol <= "D13.1 -";
10'b1011001001 : symbol <= "D13.1 +";
10'b1011000101 : symbol <= "D13.2 -";
10'b1011000101 : symbol <= "D13.2 +";
10'b1011001100 : symbol <= "D13.3 -";
10'b1011000011 : symbol <= "D13.3 +";
10'b1011001101 : symbol <= "D13.4 -";
10'b1011000010 : symbol <= "D13.4 +";
10'b1011001010 : symbol <= "D13.5 -";
10'b1011001010 : symbol <= "D13.5 +";
10'b1011000110 : symbol <= "D13.6 -";
10'b1011000110 : symbol <= "D13.6 +";
10'b1011001110 : symbol <= "D13.7 -";
10'b1011001000 : symbol <= "D13.7 +";
10'b0111001011 : symbol <= "D14.0 -";
10'b0111000100 : symbol <= "D14.0 +";
10'b0111001001 : symbol <= "D14.1 -";
10'b0111001001 : symbol <= "D14.1 +";
10'b0111000101 : symbol <= "D14.2 -";
10'b0111000101 : symbol <= "D14.2 +";
10'b0111001100 : symbol <= "D14.3 -";
10'b0111000011 : symbol <= "D14.3 +";
10'b0111001101 : symbol <= "D14.4 -";
10'b0111000010 : symbol <= "D14.4 +";
10'b0111001010 : symbol <= "D14.5 -";
10'b0111001010 : symbol <= "D14.5 +";
10'b0111000110 : symbol <= "D14.6 -";
10'b0111000110 : symbol <= "D14.6 +";
10'b0111001110 : symbol <= "D14.7 -";
10'b0111001000 : symbol <= "D14.7 +";
10'b0101110100 : symbol <= "D15.0 -";
10'b1010001011 : symbol <= "D15.0 +";
10'b0101111001 : symbol <= "D15.1 -";
10'b1010001001 : symbol <= "D15.1 +";
10'b0101110101 : symbol <= "D15.2 -";
10'b1010000101 : symbol <= "D15.2 +";
10'b0101110011 : symbol <= "D15.3 -";
10'b1010001100 : symbol <= "D15.3 +";
10'b0101110010 : symbol <= "D15.4 -";
10'b1010001101 : symbol <= "D15.4 +";
10'b0101111010 : symbol <= "D15.5 -";
10'b1010001010 : symbol <= "D15.5 +";
10'b0101110110 : symbol <= "D15.6 -";
10'b1010000110 : symbol <= "D15.6 +";
10'b0101110001 : symbol <= "D15.7 -";
10'b1010001110 : symbol <= "D15.7 +";
10'b0110110100 : symbol <= "D16.0 -";
10'b1001001011 : symbol <= "D16.0 +";
10'b0110111001 : symbol <= "D16.1 -";
10'b1001001001 : symbol <= "D16.1 +";
10'b0110110101 : symbol <= "D16.2 -";
10'b1001000101 : symbol <= "D16.2 +";
10'b0110110011 : symbol <= "D16.3 -";
10'b1001001100 : symbol <= "D16.3 +";
10'b0110110010 : symbol <= "D16.4 -";
10'b1001001101 : symbol <= "D16.4 +";
10'b0110111010 : symbol <= "D16.5 -";
10'b1001001010 : symbol <= "D16.5 +";
10'b0110110110 : symbol <= "D16.6 -";
10'b1001000110 : symbol <= "D16.6 +";
10'b0110110001 : symbol <= "D16.7 -";
10'b1001001110 : symbol <= "D16.7 +";
10'b1000111011 : symbol <= "D17.0 -";
10'b1000110100 : symbol <= "D17.0 +";
10'b1000111001 : symbol <= "D17.1 -";
10'b1000111001 : symbol <= "D17.1 +";
10'b1000110101 : symbol <= "D17.2 -";
10'b1000110101 : symbol <= "D17.2 +";
10'b1000111100 : symbol <= "D17.3 -";
10'b1000110011 : symbol <= "D17.3 +";
10'b1000111101 : symbol <= "D17.4 -";
10'b1000110010 : symbol <= "D17.4 +";
10'b1000111010 : symbol <= "D17.5 -";
10'b1000111010 : symbol <= "D17.5 +";
10'b1000110110 : symbol <= "D17.6 -";
10'b1000110110 : symbol <= "D17.6 +";
10'b1000110111 : symbol <= "D17.7 -";
10'b1000110001 : symbol <= "D17.7 +";
10'b0100111011 : symbol <= "D18.0 -";
10'b0100110100 : symbol <= "D18.0 +";
10'b0100111001 : symbol <= "D18.1 -";
10'b0100111001 : symbol <= "D18.1 +";
10'b0100110101 : symbol <= "D18.2 -";
10'b0100110101 : symbol <= "D18.2 +";
10'b0100111100 : symbol <= "D18.3 -";
10'b0100110011 : symbol <= "D18.3 +";
10'b0100111101 : symbol <= "D18.4 -";
10'b0100110010 : symbol <= "D18.4 +";
10'b0100111010 : symbol <= "D18.5 -";
10'b0100111010 : symbol <= "D18.5 +";
10'b0100110110 : symbol <= "D18.6 -";
10'b0100110110 : symbol <= "D18.6 +";
10'b0100110111 : symbol <= "D18.7 -";
10'b0100110001 : symbol <= "D18.7 +";
10'b1100101011 : symbol <= "D19.0 -";
10'b1100100100 : symbol <= "D19.0 +";
10'b1100101001 : symbol <= "D19.1 -";
10'b1100101001 : symbol <= "D19.1 +";
10'b1100100101 : symbol <= "D19.2 -";
10'b1100100101 : symbol <= "D19.2 +";
10'b1100101100 : symbol <= "D19.3 -";
10'b1100100011 : symbol <= "D19.3 +";
10'b1100101101 : symbol <= "D19.4 -";
10'b1100100010 : symbol <= "D19.4 +";
10'b1100101010 : symbol <= "D19.5 -";
10'b1100101010 : symbol <= "D19.5 +";
10'b1100100110 : symbol <= "D19.6 -";
10'b1100100110 : symbol <= "D19.6 +";
10'b1100101110 : symbol <= "D19.7 -";
10'b1100100001 : symbol <= "D19.7 +";
10'b0010111011 : symbol <= "D20.0 -";
10'b0010110100 : symbol <= "D20.0 +";
10'b0010111001 : symbol <= "D20.1 -";
10'b0010111001 : symbol <= "D20.1 +";
10'b0010110101 : symbol <= "D20.2 -";
10'b0010110101 : symbol <= "D20.2 +";
10'b0010111100 : symbol <= "D20.3 -";
10'b0010110011 : symbol <= "D20.3 +";
10'b0010111101 : symbol <= "D20.4 -";
10'b0010110010 : symbol <= "D20.4 +";
10'b0010111010 : symbol <= "D20.5 -";
10'b0010111010 : symbol <= "D20.5 +";
10'b0010110110 : symbol <= "D20.6 -";
10'b0010110110 : symbol <= "D20.6 +";
10'b0010110111 : symbol <= "D20.7 -";
10'b0010110001 : symbol <= "D20.7 +";
10'b1010101011 : symbol <= "D21.0 -";
10'b1010100100 : symbol <= "D21.0 +";
10'b1010101001 : symbol <= "D21.1 -";
10'b1010101001 : symbol <= "D21.1 +";
10'b1010100101 : symbol <= "D21.2 -";
10'b1010100101 : symbol <= "D21.2 +";
10'b1010101100 : symbol <= "D21.3 -";
10'b1010100011 : symbol <= "D21.3 +";
10'b1010101101 : symbol <= "D21.4 -";
10'b1010100010 : symbol <= "D21.4 +";
10'b1010101010 : symbol <= "D21.5 -";
10'b1010101010 : symbol <= "D21.5 +";
10'b1010100110 : symbol <= "D21.6 -";
10'b1010100110 : symbol <= "D21.6 +";
10'b1010101110 : symbol <= "D21.7 -";
10'b1010100001 : symbol <= "D21.7 +";
10'b0110101011 : symbol <= "D22.0 -";
10'b0110100100 : symbol <= "D22.0 +";
10'b0110101001 : symbol <= "D22.1 -";
10'b0110101001 : symbol <= "D22.1 +";
10'b0110100101 : symbol <= "D22.2 -";
10'b0110100101 : symbol <= "D22.2 +";
10'b0110101100 : symbol <= "D22.3 -";
10'b0110100011 : symbol <= "D22.3 +";
10'b0110101101 : symbol <= "D22.4 -";
10'b0110100010 : symbol <= "D22.4 +";
10'b0110101010 : symbol <= "D22.5 -";
10'b0110101010 : symbol <= "D22.5 +";
10'b0110100110 : symbol <= "D22.6 -";
10'b0110100110 : symbol <= "D22.6 +";
10'b0110101110 : symbol <= "D22.7 -";
10'b0110100001 : symbol <= "D22.7 +";
10'b1110100100 : symbol <= "D23.0 -";
10'b0001011011 : symbol <= "D23.0 +";
10'b1110101001 : symbol <= "D23.1 -";
10'b0001011001 : symbol <= "D23.1 +";
10'b1110100101 : symbol <= "D23.2 -";
10'b0001010101 : symbol <= "D23.2 +";
10'b1110100011 : symbol <= "D23.3 -";
10'b0001011100 : symbol <= "D23.3 +";
10'b1110100010 : symbol <= "D23.4 -";
10'b0001011101 : symbol <= "D23.4 +";
10'b1110101010 : symbol <= "D23.5 -";
10'b0001011010 : symbol <= "D23.5 +";
10'b1110100110 : symbol <= "D23.6 -";
10'b0001010110 : symbol <= "D23.6 +";
10'b1110100001 : symbol <= "D23.7 -";
10'b0001011110 : symbol <= "D23.7 +";
10'b1100110100 : symbol <= "D24.0 -";
10'b0011001011 : symbol <= "D24.0 +";
10'b1100111001 : symbol <= "D24.1 -";
10'b0011001001 : symbol <= "D24.1 +";
10'b1100110101 : symbol <= "D24.2 -";
10'b0011000101 : symbol <= "D24.2 +";
10'b1100110011 : symbol <= "D24.3 -";
10'b0011001100 : symbol <= "D24.3 +";
10'b1100110010 : symbol <= "D24.4 -";
10'b0011001101 : symbol <= "D24.4 +";
10'b1100111010 : symbol <= "D24.5 -";
10'b0011001010 : symbol <= "D24.5 +";
10'b1100110110 : symbol <= "D24.6 -";
10'b0011000110 : symbol <= "D24.6 +";
10'b1100110001 : symbol <= "D24.7 -";
10'b0011001110 : symbol <= "D24.7 +";
10'b1001101011 : symbol <= "D25.0 -";
10'b1001100100 : symbol <= "D25.0 +";
10'b1001101001 : symbol <= "D25.1 -";
10'b1001101001 : symbol <= "D25.1 +";
10'b1001100101 : symbol <= "D25.2 -";
10'b1001100101 : symbol <= "D25.2 +";
10'b1001101100 : symbol <= "D25.3 -";
10'b1001100011 : symbol <= "D25.3 +";
10'b1001101101 : symbol <= "D25.4 -";
10'b1001100010 : symbol <= "D25.4 +";
10'b1001101010 : symbol <= "D25.5 -";
10'b1001101010 : symbol <= "D25.5 +";
10'b1001100110 : symbol <= "D25.6 -";
10'b1001100110 : symbol <= "D25.6 +";
10'b1001101110 : symbol <= "D25.7 -";
10'b1001100001 : symbol <= "D25.7 +";
10'b0101101011 : symbol <= "D26.0 -";
10'b0101100100 : symbol <= "D26.0 +";
10'b0101101001 : symbol <= "D26.1 -";
10'b0101101001 : symbol <= "D26.1 +";
10'b0101100101 : symbol <= "D26.2 -";
10'b0101100101 : symbol <= "D26.2 +";
10'b0101101100 : symbol <= "D26.3 -";
10'b0101100011 : symbol <= "D26.3 +";
10'b0101101101 : symbol <= "D26.4 -";
10'b0101100010 : symbol <= "D26.4 +";
10'b0101101010 : symbol <= "D26.5 -";
10'b0101101010 : symbol <= "D26.5 +";
10'b0101100110 : symbol <= "D26.6 -";
10'b0101100110 : symbol <= "D26.6 +";
10'b0101101110 : symbol <= "D26.7 -";
10'b0101100001 : symbol <= "D26.7 +";
10'b1101100100 : symbol <= "D27.0 -";
10'b0010011011 : symbol <= "D27.0 +";
10'b1101101001 : symbol <= "D27.1 -";
10'b0010011001 : symbol <= "D27.1 +";
10'b1101100101 : symbol <= "D27.2 -";
10'b0010010101 : symbol <= "D27.2 +";
10'b1101100011 : symbol <= "D27.3 -";
10'b0010011100 : symbol <= "D27.3 +";
10'b1101100010 : symbol <= "D27.4 -";
10'b0010011101 : symbol <= "D27.4 +";
10'b1101101010 : symbol <= "D27.5 -";
10'b0010011010 : symbol <= "D27.5 +";
10'b1101100110 : symbol <= "D27.6 -";
10'b0010010110 : symbol <= "D27.6 +";
10'b1101100001 : symbol <= "D27.7 -";
10'b0010011110 : symbol <= "D27.7 +";
10'b0011101011 : symbol <= "D28.0 -";
10'b0011100100 : symbol <= "D28.0 +";
10'b0011101001 : symbol <= "D28.1 -";
10'b0011101001 : symbol <= "D28.1 +";
10'b0011100101 : symbol <= "D28.2 -";
10'b0011100101 : symbol <= "D28.2 +";
10'b0011101100 : symbol <= "D28.3 -";
10'b0011100011 : symbol <= "D28.3 +";
10'b0011101101 : symbol <= "D28.4 -";
10'b0011100010 : symbol <= "D28.4 +";
10'b0011101010 : symbol <= "D28.5 -";
10'b0011101010 : symbol <= "D28.5 +";
10'b0011100110 : symbol <= "D28.6 -";
10'b0011100110 : symbol <= "D28.6 +";
10'b0011101110 : symbol <= "D28.7 -";
10'b0011100001 : symbol <= "D28.7 +";
10'b1011100100 : symbol <= "D29.0 -";
10'b0100011011 : symbol <= "D29.0 +";
10'b1011101001 : symbol <= "D29.1 -";
10'b0100011001 : symbol <= "D29.1 +";
10'b1011100101 : symbol <= "D29.2 -";
10'b0100010101 : symbol <= "D29.2 +";
10'b1011100011 : symbol <= "D29.3 -";
10'b0100011100 : symbol <= "D29.3 +";
10'b1011100010 : symbol <= "D29.4 -";
10'b0100011101 : symbol <= "D29.4 +";
10'b1011101010 : symbol <= "D29.5 -";
10'b0100011010 : symbol <= "D29.5 +";
10'b1011100110 : symbol <= "D29.6 -";
10'b0100010110 : symbol <= "D29.6 +";
10'b1011100001 : symbol <= "D29.7 -";
10'b0100011110 : symbol <= "D29.7 +";
10'b0111100100 : symbol <= "D30.0 -";
10'b1000011011 : symbol <= "D30.0 +";
10'b0111101001 : symbol <= "D30.1 -";
10'b1000011001 : symbol <= "D30.1 +";
10'b0111100101 : symbol <= "D30.2 -";
10'b1000010101 : symbol <= "D30.2 +";
10'b0111100011 : symbol <= "D30.3 -";
10'b1000011100 : symbol <= "D30.3 +";
10'b0111100010 : symbol <= "D30.4 -";
10'b1000011101 : symbol <= "D30.4 +";
10'b0111101010 : symbol <= "D30.5 -";
10'b1000011010 : symbol <= "D30.5 +";
10'b0111100110 : symbol <= "D30.6 -";
10'b1000010110 : symbol <= "D30.6 +";
10'b0111100001 : symbol <= "D30.7 -";
10'b1000011110 : symbol <= "D30.7 +";
10'b1010110100 : symbol <= "D31.0 -";
10'b0101001011 : symbol <= "D31.0 +";
10'b1010111001 : symbol <= "D31.1 -";
10'b0101001001 : symbol <= "D31.1 +";
10'b1010110101 : symbol <= "D31.2 -";
10'b0101000101 : symbol <= "D31.2 +";
10'b1010110011 : symbol <= "D31.3 -";
10'b0101001100 : symbol <= "D31.3 +";
10'b1010110010 : symbol <= "D31.4 -";
10'b0101001101 : symbol <= "D31.4 +";
10'b1010111010 : symbol <= "D31.5 -";
10'b0101001010 : symbol <= "D31.5 +";
10'b1010110110 : symbol <= "D31.6 -";
10'b0101000110 : symbol <= "D31.6 +";
10'b1010110001 : symbol <= "D31.7 -";
10'b0101001110 : symbol <= "D31.7 +";
10'b0011110100 : symbol <= "K28.0 -";
10'b0011111001 : symbol <= "K28.1 -";
10'b0011110101 : symbol <= "K28.2 -";
10'b0011110011 : symbol <= "K28.3 -";
10'b0011110010 : symbol <= "K28.4 -";
10'b0011111010 : symbol <= "K28.5 -";
10'b0011110110 : symbol <= "K28.6 -";
10'b0011111000 : symbol <= "K28.7 -";
10'b1110101000 : symbol <= "K23.7 -";
10'b1101101000 : symbol <= "K27.7 -";
10'b1011101000 : symbol <= "K29.7 -";
10'b0111101000 : symbol <= "K30.7 -";
10'b1100001011 : symbol <= "K28.0 +";
10'b1100000110 : symbol <= "K28.1 +";
10'b1100001010 : symbol <= "K28.2 +";
10'b1100001100 : symbol <= "K28.3 +";
10'b1100001101 : symbol <= "K28.4 +";
10'b1100000101 : symbol <= "K28.5 +";
10'b1100001001 : symbol <= "K28.6 +";
10'b1100000111 : symbol <= "K28.7 +";
10'b0001010111 : symbol <= "K23.7 +";
10'b0010010111 : symbol <= "K27.7 +";
10'b0100010111 : symbol <= "K29.7 +";
10'b1000010111 : symbol <= "K30.7 +";
